// Copyright (C) 2023  Intel Corporation. All rights reserved.
// Your use of Intel Corporation's design tools, logic functions 
// and other software and tools, and any partner logic 
// functions, and any output files from any of the foregoing 
// (including device programming or simulation files), and any 
// associated documentation or information are expressly subject 
// to the terms and conditions of the Intel Program License 
// Subscription Agreement, the Intel Quartus Prime License Agreement,
// the Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is for
// the sole purpose of programming logic devices manufactured by
// Intel and sold by Intel or its authorized distributors.  Please
// refer to the applicable agreement for further details, at
// https://fpgasoftware.intel.com/eula.

// PROGRAM		"Quartus Prime"
// VERSION		"Version 22.1std.1 Build 917 02/14/2023 SC Lite Edition"
// CREATED		"Thu Mar 30 19:43:44 2023"

module ALU_74181(
	S3,
	S2,
	S1,
	S0,
	B3N,
	A3N,
	B2N,
	A2N,
	B1N,
	A1N,
	B0N,
	A0N,
	CN,
	M,
	F1N,
	AEQB,
	F2N,
	F3N,
	PN,
	CN4,
	GN,
	F0N
);


input wire	S3;
input wire	S2;
input wire	S1;
input wire	S0;
input wire	B3N;
input wire	A3N;
input wire	B2N;
input wire	A2N;
input wire	B1N;
input wire	A1N;
input wire	B0N;
input wire	A0N;
input wire	CN;
input wire	M;
output wire	F1N;
output wire	AEQB;
output wire	F2N;
output wire	F3N;
output wire	PN;
output wire	CN4;
output wire	GN;
output wire	F0N;

wire	SYNTHESIZED_WIRE_117;
wire	SYNTHESIZED_WIRE_118;
wire	SYNTHESIZED_WIRE_119;
wire	SYNTHESIZED_WIRE_6;
wire	SYNTHESIZED_WIRE_7;
wire	SYNTHESIZED_WIRE_8;
wire	SYNTHESIZED_WIRE_9;
wire	SYNTHESIZED_WIRE_10;
wire	SYNTHESIZED_WIRE_11;
wire	SYNTHESIZED_WIRE_12;
wire	SYNTHESIZED_WIRE_13;
wire	SYNTHESIZED_WIRE_14;
wire	SYNTHESIZED_WIRE_15;
wire	SYNTHESIZED_WIRE_16;
wire	SYNTHESIZED_WIRE_17;
wire	SYNTHESIZED_WIRE_18;
wire	SYNTHESIZED_WIRE_19;
wire	SYNTHESIZED_WIRE_20;
wire	SYNTHESIZED_WIRE_21;
wire	SYNTHESIZED_WIRE_22;
wire	SYNTHESIZED_WIRE_23;
wire	SYNTHESIZED_WIRE_24;
wire	SYNTHESIZED_WIRE_25;
wire	SYNTHESIZED_WIRE_26;
wire	SYNTHESIZED_WIRE_27;
wire	SYNTHESIZED_WIRE_28;
wire	SYNTHESIZED_WIRE_29;
wire	SYNTHESIZED_WIRE_120;
wire	SYNTHESIZED_WIRE_121;
wire	SYNTHESIZED_WIRE_122;
wire	SYNTHESIZED_WIRE_123;
wire	SYNTHESIZED_WIRE_124;
wire	SYNTHESIZED_WIRE_125;
wire	SYNTHESIZED_WIRE_126;
wire	SYNTHESIZED_WIRE_127;
wire	SYNTHESIZED_WIRE_56;
wire	SYNTHESIZED_WIRE_57;
wire	SYNTHESIZED_WIRE_58;
wire	SYNTHESIZED_WIRE_128;
wire	SYNTHESIZED_WIRE_129;
wire	SYNTHESIZED_WIRE_86;
wire	SYNTHESIZED_WIRE_87;
wire	SYNTHESIZED_WIRE_88;
wire	SYNTHESIZED_WIRE_89;
wire	SYNTHESIZED_WIRE_90;
wire	SYNTHESIZED_WIRE_91;
wire	SYNTHESIZED_WIRE_92;
wire	SYNTHESIZED_WIRE_93;
wire	SYNTHESIZED_WIRE_94;
wire	SYNTHESIZED_WIRE_95;
wire	SYNTHESIZED_WIRE_96;
wire	SYNTHESIZED_WIRE_97;
wire	SYNTHESIZED_WIRE_98;
wire	SYNTHESIZED_WIRE_99;
wire	SYNTHESIZED_WIRE_101;
wire	SYNTHESIZED_WIRE_102;
wire	SYNTHESIZED_WIRE_103;
wire	SYNTHESIZED_WIRE_104;
wire	SYNTHESIZED_WIRE_105;
wire	SYNTHESIZED_WIRE_106;
wire	SYNTHESIZED_WIRE_107;
wire	SYNTHESIZED_WIRE_108;
wire	SYNTHESIZED_WIRE_109;
wire	SYNTHESIZED_WIRE_110;
wire	SYNTHESIZED_WIRE_111;
wire	SYNTHESIZED_WIRE_112;
wire	SYNTHESIZED_WIRE_113;
wire	SYNTHESIZED_WIRE_114;
wire	SYNTHESIZED_WIRE_115;
wire	SYNTHESIZED_WIRE_116;

assign	F1N = SYNTHESIZED_WIRE_109;
assign	F2N = SYNTHESIZED_WIRE_108;
assign	F3N = SYNTHESIZED_WIRE_107;
assign	GN = SYNTHESIZED_WIRE_96;
assign	F0N = SYNTHESIZED_WIRE_110;



assign	SYNTHESIZED_WIRE_14 = S0 & B1N;

assign	SYNTHESIZED_WIRE_15 = SYNTHESIZED_WIRE_117 & S1;

assign	SYNTHESIZED_WIRE_21 = SYNTHESIZED_WIRE_117 & S2 & A1N;

assign	SYNTHESIZED_WIRE_20 = A1N & S3 & B1N;

assign	SYNTHESIZED_WIRE_16 = S0 & B2N;

assign	SYNTHESIZED_WIRE_17 = SYNTHESIZED_WIRE_118 & S1;

assign	SYNTHESIZED_WIRE_23 = SYNTHESIZED_WIRE_118 & S2 & A2N;

assign	SYNTHESIZED_WIRE_22 = A2N & S3 & B2N;

assign	SYNTHESIZED_WIRE_26 = S0 & B3N;

assign	SYNTHESIZED_WIRE_27 = SYNTHESIZED_WIRE_119 & S1;

assign	SYNTHESIZED_WIRE_29 = SYNTHESIZED_WIRE_119 & S2 & A3N;

assign	SYNTHESIZED_WIRE_28 = A3N & S3 & B3N;

assign	SYNTHESIZED_WIRE_119 =  ~B3N;

assign	SYNTHESIZED_WIRE_129 =  ~B0N;

assign	SYNTHESIZED_WIRE_117 =  ~B1N;

assign	SYNTHESIZED_WIRE_118 =  ~B2N;


soft	b2v_37(
	.in(SYNTHESIZED_WIRE_6),
	.out(SYNTHESIZED_WIRE_121));


soft	b2v_38(
	.in(SYNTHESIZED_WIRE_7),
	.out(SYNTHESIZED_WIRE_120));


soft	b2v_39(
	.in(SYNTHESIZED_WIRE_8),
	.out(SYNTHESIZED_WIRE_123));


soft	b2v_40(
	.in(SYNTHESIZED_WIRE_9),
	.out(SYNTHESIZED_WIRE_122));


soft	b2v_41(
	.in(SYNTHESIZED_WIRE_10),
	.out(SYNTHESIZED_WIRE_125));


soft	b2v_42(
	.in(SYNTHESIZED_WIRE_11),
	.out(SYNTHESIZED_WIRE_124));

assign	SYNTHESIZED_WIRE_6 = ~(A0N | SYNTHESIZED_WIRE_12 | SYNTHESIZED_WIRE_13);

assign	SYNTHESIZED_WIRE_8 = ~(A1N | SYNTHESIZED_WIRE_14 | SYNTHESIZED_WIRE_15);

assign	SYNTHESIZED_WIRE_10 = ~(A2N | SYNTHESIZED_WIRE_16 | SYNTHESIZED_WIRE_17);

assign	SYNTHESIZED_WIRE_7 = ~(SYNTHESIZED_WIRE_18 | SYNTHESIZED_WIRE_19);

assign	SYNTHESIZED_WIRE_9 = ~(SYNTHESIZED_WIRE_20 | SYNTHESIZED_WIRE_21);

assign	SYNTHESIZED_WIRE_11 = ~(SYNTHESIZED_WIRE_22 | SYNTHESIZED_WIRE_23);


soft	b2v_49(
	.in(SYNTHESIZED_WIRE_24),
	.out(SYNTHESIZED_WIRE_126));


soft	b2v_50(
	.in(SYNTHESIZED_WIRE_25),
	.out(SYNTHESIZED_WIRE_127));

assign	SYNTHESIZED_WIRE_25 = ~(A3N | SYNTHESIZED_WIRE_26 | SYNTHESIZED_WIRE_27);

assign	SYNTHESIZED_WIRE_24 = ~(SYNTHESIZED_WIRE_28 | SYNTHESIZED_WIRE_29);

assign	SYNTHESIZED_WIRE_101 = SYNTHESIZED_WIRE_120 ^ SYNTHESIZED_WIRE_121;

assign	SYNTHESIZED_WIRE_103 = SYNTHESIZED_WIRE_122 ^ SYNTHESIZED_WIRE_123;

assign	SYNTHESIZED_WIRE_105 = SYNTHESIZED_WIRE_124 ^ SYNTHESIZED_WIRE_125;

assign	SYNTHESIZED_WIRE_94 = SYNTHESIZED_WIRE_126 ^ SYNTHESIZED_WIRE_127;

assign	SYNTHESIZED_WIRE_56 = SYNTHESIZED_WIRE_126 & SYNTHESIZED_WIRE_125;

assign	SYNTHESIZED_WIRE_57 = SYNTHESIZED_WIRE_123 & SYNTHESIZED_WIRE_124 & SYNTHESIZED_WIRE_126;

assign	SYNTHESIZED_WIRE_12 = S0 & B0N;

assign	PN = ~(SYNTHESIZED_WIRE_126 & SYNTHESIZED_WIRE_124 & SYNTHESIZED_WIRE_122 & SYNTHESIZED_WIRE_120);

assign	SYNTHESIZED_WIRE_97 = ~(SYNTHESIZED_WIRE_124 & SYNTHESIZED_WIRE_122 & SYNTHESIZED_WIRE_120 & SYNTHESIZED_WIRE_126 & CN & CN);

assign	SYNTHESIZED_WIRE_58 = SYNTHESIZED_WIRE_126 & SYNTHESIZED_WIRE_124 & SYNTHESIZED_WIRE_122 & SYNTHESIZED_WIRE_121;

assign	SYNTHESIZED_WIRE_96 = ~(SYNTHESIZED_WIRE_127 | SYNTHESIZED_WIRE_56 | SYNTHESIZED_WIRE_57 | SYNTHESIZED_WIRE_58);

assign	SYNTHESIZED_WIRE_102 = ~(CN & SYNTHESIZED_WIRE_128);

assign	SYNTHESIZED_WIRE_99 = SYNTHESIZED_WIRE_121 & SYNTHESIZED_WIRE_128;

assign	SYNTHESIZED_WIRE_98 = SYNTHESIZED_WIRE_128 & SYNTHESIZED_WIRE_120 & CN;

assign	SYNTHESIZED_WIRE_90 = SYNTHESIZED_WIRE_123 & SYNTHESIZED_WIRE_128;

assign	SYNTHESIZED_WIRE_91 = SYNTHESIZED_WIRE_128 & SYNTHESIZED_WIRE_121 & SYNTHESIZED_WIRE_122;

assign	SYNTHESIZED_WIRE_92 = CN & SYNTHESIZED_WIRE_120 & SYNTHESIZED_WIRE_122 & SYNTHESIZED_WIRE_128;

assign	SYNTHESIZED_WIRE_13 = SYNTHESIZED_WIRE_129 & S1;

assign	SYNTHESIZED_WIRE_89 = SYNTHESIZED_WIRE_125 & SYNTHESIZED_WIRE_128;

assign	SYNTHESIZED_WIRE_88 = SYNTHESIZED_WIRE_128 & SYNTHESIZED_WIRE_123 & SYNTHESIZED_WIRE_124;

assign	SYNTHESIZED_WIRE_87 = SYNTHESIZED_WIRE_122 & SYNTHESIZED_WIRE_124 & SYNTHESIZED_WIRE_121 & SYNTHESIZED_WIRE_128;

assign	SYNTHESIZED_WIRE_86 = CN & SYNTHESIZED_WIRE_120 & SYNTHESIZED_WIRE_122 & CN & SYNTHESIZED_WIRE_124 & SYNTHESIZED_WIRE_128;

assign	SYNTHESIZED_WIRE_93 = ~(SYNTHESIZED_WIRE_86 | SYNTHESIZED_WIRE_87 | SYNTHESIZED_WIRE_88 | SYNTHESIZED_WIRE_89);

assign	SYNTHESIZED_WIRE_116 = ~(SYNTHESIZED_WIRE_90 | SYNTHESIZED_WIRE_91 | SYNTHESIZED_WIRE_92);


soft	b2v_76(
	.in(SYNTHESIZED_WIRE_93),
	.out(SYNTHESIZED_WIRE_95));

assign	SYNTHESIZED_WIRE_111 = SYNTHESIZED_WIRE_94 ^ SYNTHESIZED_WIRE_95;

assign	CN4 = ~(SYNTHESIZED_WIRE_96 & SYNTHESIZED_WIRE_97);

assign	SYNTHESIZED_WIRE_115 = ~(SYNTHESIZED_WIRE_98 | SYNTHESIZED_WIRE_99);

assign	SYNTHESIZED_WIRE_19 = SYNTHESIZED_WIRE_129 & S2 & A0N;

assign	SYNTHESIZED_WIRE_114 = SYNTHESIZED_WIRE_101 ^ SYNTHESIZED_WIRE_102;

assign	SYNTHESIZED_WIRE_113 = SYNTHESIZED_WIRE_103 ^ SYNTHESIZED_WIRE_104;

assign	SYNTHESIZED_WIRE_112 = SYNTHESIZED_WIRE_105 ^ SYNTHESIZED_WIRE_106;

assign	AEQB = SYNTHESIZED_WIRE_107 & SYNTHESIZED_WIRE_108 & SYNTHESIZED_WIRE_109 & SYNTHESIZED_WIRE_110;


soft	b2v_84(
	.in(SYNTHESIZED_WIRE_111),
	.out(SYNTHESIZED_WIRE_107));


soft	b2v_85(
	.in(SYNTHESIZED_WIRE_112),
	.out(SYNTHESIZED_WIRE_108));


soft	b2v_86(
	.in(SYNTHESIZED_WIRE_113),
	.out(SYNTHESIZED_WIRE_109));


soft	b2v_87(
	.in(SYNTHESIZED_WIRE_114),
	.out(SYNTHESIZED_WIRE_110));


soft	b2v_88(
	.in(SYNTHESIZED_WIRE_115),
	.out(SYNTHESIZED_WIRE_104));


soft	b2v_89(
	.in(SYNTHESIZED_WIRE_116),
	.out(SYNTHESIZED_WIRE_106));

assign	SYNTHESIZED_WIRE_18 = A0N & S3 & B0N;

assign	SYNTHESIZED_WIRE_128 =  ~M;


endmodule